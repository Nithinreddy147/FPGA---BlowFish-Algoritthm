`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.04.2024 01:12:51
// Design Name: 
// Module Name: BLFH
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// Module for key expansion
module blowfish_key_expansion (
    input [31:0] key,         // Input key
    output reg [31:0] subkeys // Generated subkeys
);
    reg [31:0] P [17:0];  // P-array
    reg [31:0] temp;
    integer i;
    
    // Initial P-array values
    initial begin
        P[0]  = 32'h243f6a88;
        P[1]  = 32'h85a308d3;
        P[2]  = 32'h13198a2e;
        P[3]  = 32'h03707344;
        P[4]  = 32'ha4093822;
        P[5]  = 32'h299f31d0;
        P[6]  = 32'h082efa98;
        P[7]  = 32'hec4e6c89;
        P[8]  = 32'h452821e6;
        P[9]  = 32'h38d01377;
        P[10] = 32'hbe5466cf;
        P[11] = 32'h34e90c6c;
        P[12] = 32'hc0ac29b7;
        P[13] = 32'hc97c50dd;
        P[14] = 32'h3f84d5b5;
        P[15] = 32'hb5470917;
        P[16] = 32'h9216d5d9;
        P[17] = 32'h8979fb1b;
    end

    // Key schedule algorithm
    always @(*) begin
        // Initialize P-array with initial values
        for (i = 0; i < 18; i = i + 1) begin
            P[i] = P[i] ^ key[(i*32) +: 32];
        end
        
        // Expand key into subkeys
        temp = 32'h0;
        for (i = 0; i < 18; i = i + 1) begin
            temp = temp ^ P[i];
            subkeys[i] = temp;
        end
    end
endmodule

// Module for Blowfish encryption
module blowfish_encrypt(
    input [63:0] plaintext,               // Input plaintext
    input [31:0] subkeys [17:0],          // Subkeys generated by key expansion
    output reg [63:0] ciphertext          // Output ciphertext
);
    reg [31:0] L, R;
    integer i;
    
    // Declare S-box arrays
    reg [31:0] S0 [255:0];
    reg [31:0] S1 [255:0];
    reg [31:0] S2 [255:0];
    reg [31:0] S3 [255:0];
    
    // Initial permutation
    initial begin
        L = plaintext[63:32];
        R = plaintext[31:0];
    end
    
    // Read S-box values from text file and initialize S-box arrays
    initial begin
        $readmemh("sbox1.txt", S0);
        $readmemh("sbox2.txt", S1);
        $readmemh("sbox3.txt", S2);
        $readmemh("sbox4.txt", S3);
    end

    // 16 rounds of encryption
    always @(*) begin
        for (i = 0; i < 16; i = i + 1) begin
            L = L ^ subkeys[i];
            R = R ^ F(L);
            {L, R} = {R, L}; // Swap L and R
        end
        {L, R} = {R, L}; // Swap L and R back after the last round
        L = L ^ subkeys[16];
        R = R ^ subkeys[17];
        ciphertext = {L, R};
    end

    // Function for the F function
    function [31:0] F;
    input [31:0] x;
    reg [7:0] b0, b1, b2, b3;
    reg [7:0] sb0, sb1, sb2, sb3;
    reg [31:0] result;
    begin
        // Split the 32-bit input into four 8-bit segments
        b0 = x[31:24];
        b1 = x[23:16];
        b2 = x[15:8];
        b3 = x[7:0];

        // Apply the four S-boxes to each 8-bit segment
        sb0 = S0[b0];
        sb1 = S1[b1];
        sb2 = S2[b2];
        sb3 = S3[b3];

        // Combine the results from the S-boxes
        result = {sb0, sb1, sb2, sb3};

        // Apply a permutation to the result
        result = permutation(result);

        F = result;
    end
    endfunction
    
    // Function for permutation using the P-array
    function [31:0] permutation;
        input [31:0] x;
        reg [7:0] b0, b1, b2, b3;
        reg [7:0] sb0, sb1, sb2, sb3;
        reg [31:0] result;
        begin
            // Split the 32-bit input into four 8-bit segments
            b0 = x[31:24];
            b1 = x[23:16];
            b2 = x[15:8];
            b3 = x[7:0];
    
            // Apply the four S-boxes to each 8-bit segment
            sb0 = S0[b0];
            sb1 = S1[b1];
            sb2 = S2[b2];
            sb3 = S3[b3];
    
            // Combine the results from the S-boxes
            result = {sb0, sb1, sb2, sb3};
    
            // Apply a permutation to the result
            result = {
            result[7:0],     // Take the least significant byte of the result
            result[15:8],    // Take the third least significant byte of the result
            result[23:16],   // Take the second least significant byte of the result
            result[31:24]    // Take the most significant byte of the result
        };
    
            permutation = result;
        end
    endfunction
endmodule

// Module for Blowfish decryption
module blowfish_decrypt(
    input [63:0] ciphertext,               // Input ciphertext
    input [31:0] subkeys [17:0],           // Subkeys generated by key expansion (in reverse order)
    output reg [63:0] plaintext            // Output plaintext
);
    reg [31:0] L, R;
    integer i;
    
    // Declare S-box arrays (same as in encryption module)
    reg [31:0] S0 [255:0];
    reg [31:0] S1 [255:0];
    reg [31:0] S2 [255:0];
    reg [31:0] S3 [255:0];
    
    // Initial permutation (same as in encryption module)
    initial begin
        L = ciphertext[63:32];
        R = ciphertext[31:0];
    end
    
    // Read S-box values from text file and initialize S-box arrays (same as in encryption module)
    initial begin
        $readmemh("sbox1.txt", S0);
        $readmemh("sbox2.txt", S1);
        $readmemh("sbox3.txt", S2);
        $readmemh("sbox4.txt", S3);
    end

    // 16 rounds of decryption (same as in encryption module, but with subkeys used in reverse order)
    always @(*) begin
        for (i = 17; i > 1; i = i - 1) begin
            L = L ^ subkeys[i];
            R = R ^ F(L);
            {L, R} = {R, L}; // Swap L and R
        end
        {L, R} = {R, L}; // Swap L and R back after the last round
        L = L ^ subkeys[1];
        R = R ^ subkeys[0];
        plaintext = {L, R};
    end

    // Function for the F function (same as in encryption module)
    function [31:0] F;
    input [31:0] x;
    reg [7:0] b0, b1, b2, b3;
    reg [7:0] sb0, sb1, sb2, sb3;
    reg [31:0] result;
    begin
        // Split the 32-bit input into four 8-bit segments
        b0 = x[31:24];
        b1 = x[23:16];
        b2 = x[15:8];
        b3 = x[7:0];

        // Apply the four S-boxes to each 8-bit segment
        sb0 = S0[b0];
        sb1 = S1[b1];
        sb2 = S2[b2];
        sb3 = S3[b3];

        // Combine the results from the S-boxes
        result = {sb0, sb1, sb2, sb3};

        // Apply a permutation to the result (same as in encryption module)
        result = {
            result[7:0],    // Take the least significant byte of the result
            result[15:8],   // Take the third least significant byte of the result
            result[23:16],  // Take the second least significant byte of the result
            result[31:24]   // Take the most significant byte of the result
        };

        F = result;
    end
    endfunction
endmodule

